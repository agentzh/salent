library verilog;
use verilog.vl_types.all;
entity read_byte is
end read_byte;
