library verilog;
use verilog.vl_types.all;
entity idu is
    generic(
        addr_size       : integer := 32;
        \DISP_LEN\      : integer := 4;
        \IMM_LEN\       : integer := 6;
        syntax_error    : integer := 0;
        end_error       : integer := 1;
        s_0             : integer := 0;
        s_1             : integer := 1;
        s_2             : integer := 2;
        s_3             : integer := 3;
        s_4             : integer := 4;
        s_5             : integer := 5;
        s_6             : integer := 6;
        s_7             : integer := 7;
        s_8             : integer := 8;
        s_9             : integer := 9;
        s_10            : integer := 10;
        s_11            : integer := 11;
        s_12            : integer := 12;
        s_13            : integer := 13;
        s_14            : integer := 14;
        s_15            : integer := 15;
        s_16            : integer := 16;
        s_17            : integer := 17;
        s_18            : integer := 18;
        s_19            : integer := 19;
        s_20            : integer := 20;
        s_21            : integer := 21;
        s_22            : integer := 22;
        s_23            : integer := 23;
        s_24            : integer := 24;
        s_25            : integer := 25;
        s_26            : integer := 26;
        s_27            : integer := 27;
        s_28            : integer := 28;
        s_29            : integer := 29;
        s_30            : integer := 30;
        s_31            : integer := 31;
        s_32            : integer := 32;
        s_33            : integer := 33;
        s_34            : integer := 34;
        s_35            : integer := 35;
        s_36            : integer := 36;
        s_37            : integer := 37;
        s_38            : integer := 38;
        s_39            : integer := 39;
        s_40            : integer := 40;
        s_41            : integer := 41;
        s_42            : integer := 42;
        s_43            : integer := 43;
        s_44            : integer := 44;
        s_45            : integer := 45;
        s_46            : integer := 46;
        s_47            : integer := 47;
        s_48            : integer := 48;
        s_49            : integer := 49;
        s_50            : integer := 50;
        s_51            : integer := 51;
        s_52            : integer := 52;
        s_53            : integer := 53;
        s_54            : integer := 54;
        s_55            : integer := 55;
        s_56            : integer := 56;
        s_57            : integer := 57;
        s_58            : integer := 58;
        s_59            : integer := 59;
        s_60            : integer := 60;
        s_61            : integer := 61;
        s_62            : integer := 62;
        s_63            : integer := 63;
        s_64            : integer := 64;
        s_65            : integer := 65;
        s_66            : integer := 66;
        s_67            : integer := 67;
        s_68            : integer := 68;
        s_69            : integer := 69;
        s_70            : integer := 70;
        s_71            : integer := 71;
        s_72            : integer := 72;
        s_73            : integer := 73;
        s_74            : integer := 74;
        s_75            : integer := 75;
        s_76            : integer := 76;
        s_77            : integer := 77;
        s_78            : integer := 78;
        s_79            : integer := 79;
        s_80            : integer := 80;
        s_81            : integer := 81;
        s_82            : integer := 82;
        s_83            : integer := 83;
        s_84            : integer := 84;
        s_85            : integer := 85;
        s_86            : integer := 86;
        s_87            : integer := 87;
        s_88            : integer := 88;
        s_89            : integer := 89;
        s_90            : integer := 90;
        s_91            : integer := 91;
        s_92            : integer := 92;
        s_93            : integer := 93;
        s_94            : integer := 94;
        s_95            : integer := 95;
        s_96            : integer := 96;
        s_97            : integer := 97;
        s_98            : integer := 98;
        s_99            : integer := 99;
        s_100           : integer := 100;
        s_101           : integer := 101;
        s_102           : integer := 102;
        s_103           : integer := 103;
        s_104           : integer := 104;
        s_105           : integer := 105;
        s_106           : integer := 106;
        s_107           : integer := 107;
        s_108           : integer := 108;
        s_109           : integer := 109;
        s_110           : integer := 110;
        s_111           : integer := 111;
        s_112           : integer := 112;
        s_113           : integer := 113;
        s_114           : integer := 114;
        s_115           : integer := 115;
        s_116           : integer := 116;
        s_117           : integer := 117;
        s_118           : integer := 118;
        s_119           : integer := 119;
        s_120           : integer := 120;
        s_121           : integer := 121;
        s_122           : integer := 122;
        s_123           : integer := 123;
        s_124           : integer := 124;
        s_125           : integer := 125;
        s_126           : integer := 126;
        s_127           : integer := 127;
        s_128           : integer := 128;
        s_129           : integer := 129;
        s_130           : integer := 130;
        s_131           : integer := 131;
        s_132           : integer := 132;
        s_133           : integer := 133;
        s_134           : integer := 134;
        s_135           : integer := 135;
        s_136           : integer := 136;
        s_137           : integer := 137;
        s_138           : integer := 138;
        s_139           : integer := 139;
        s_140           : integer := 140;
        s_141           : integer := 141;
        s_142           : integer := 142;
        s_143           : integer := 143;
        s_144           : integer := 144;
        s_145           : integer := 145;
        s_146           : integer := 146;
        s_147           : integer := 147;
        s_148           : integer := 148;
        s_149           : integer := 149;
        s_150           : integer := 150;
        s_151           : integer := 151;
        s_152           : integer := 152;
        s_153           : integer := 153;
        s_154           : integer := 154;
        s_155           : integer := 155;
        s_156           : integer := 156;
        s_157           : integer := 157;
        s_158           : integer := 158;
        s_159           : integer := 159;
        s_160           : integer := 160;
        s_161           : integer := 161;
        s_162           : integer := 162;
        s_163           : integer := 163;
        s_164           : integer := 164;
        s_165           : integer := 165;
        s_166           : integer := 166;
        s_167           : integer := 167;
        s_168           : integer := 168;
        s_169           : integer := 169;
        s_170           : integer := 170;
        s_171           : integer := 171;
        s_172           : integer := 172;
        s_173           : integer := 173;
        s_174           : integer := 174;
        s_175           : integer := 175;
        s_176           : integer := 176;
        s_177           : integer := 177;
        s_178           : integer := 178;
        s_179           : integer := 179;
        s_180           : integer := 180;
        s_181           : integer := 181;
        s_182           : integer := 182;
        s_183           : integer := 183;
        s_184           : integer := 184;
        s_185           : integer := 185;
        s_186           : integer := 186;
        s_187           : integer := 187;
        s_188           : integer := 188;
        s_189           : integer := 189;
        s_190           : integer := 190;
        s_191           : integer := 191;
        s_192           : integer := 192;
        s_193           : integer := 193;
        s_194           : integer := 194;
        s_195           : integer := 195;
        s_196           : integer := 196;
        s_197           : integer := 197;
        s_198           : integer := 198;
        s_199           : integer := 199;
        s_200           : integer := 200;
        s_201           : integer := 201;
        s_202           : integer := 202;
        s_203           : integer := 203;
        s_204           : integer := 204;
        s_205           : integer := 205;
        s_206           : integer := 206;
        s_207           : integer := 207;
        s_208           : integer := 208;
        s_209           : integer := 209;
        s_210           : integer := 210;
        s_211           : integer := 211;
        s_212           : integer := 212;
        s_213           : integer := 213;
        s_214           : integer := 214;
        s_215           : integer := 215;
        s_216           : integer := 216;
        s_217           : integer := 217;
        s_218           : integer := 218;
        s_219           : integer := 219;
        s_220           : integer := 220;
        s_221           : integer := 221;
        s_222           : integer := 222;
        s_223           : integer := 223;
        s_224           : integer := 224;
        s_225           : integer := 225;
        s_226           : integer := 226;
        s_227           : integer := 227;
        s_228           : integer := 228;
        s_229           : integer := 229;
        s_230           : integer := 230;
        s_231           : integer := 231;
        s_232           : integer := 232;
        s_233           : integer := 233;
        s_234           : integer := 234;
        s_235           : integer := 235;
        s_236           : integer := 236;
        s_237           : integer := 237;
        s_238           : integer := 238;
        s_239           : integer := 239;
        s_240           : integer := 240;
        s_241           : integer := 241;
        s_242           : integer := 242;
        s_243           : integer := 243;
        s_244           : integer := 244;
        s_245           : integer := 245;
        s_246           : integer := 246;
        s_247           : integer := 247;
        s_248           : integer := 248;
        s_249           : integer := 249;
        s_250           : integer := 250;
        s_251           : integer := 251;
        s_252           : integer := 252;
        s_253           : integer := 253;
        s_254           : integer := 254;
        s_255           : integer := 255;
        s_256           : integer := 256;
        s_257           : integer := 257;
        s_258           : integer := 258;
        s_259           : integer := 259;
        s_260           : integer := 260;
        s_261           : integer := 261;
        s_262           : integer := 262;
        s_263           : integer := 263;
        s_264           : integer := 264;
        s_265           : integer := 265;
        s_266           : integer := 266;
        s_267           : integer := 267;
        s_268           : integer := 268;
        s_269           : integer := 269;
        s_270           : integer := 270;
        s_271           : integer := 271;
        s_272           : integer := 272;
        s_273           : integer := 273;
        s_274           : integer := 274;
        s_275           : integer := 275;
        s_276           : integer := 276;
        s_277           : integer := 277;
        s_278           : integer := 278;
        s_279           : integer := 279;
        s_280           : integer := 280;
        s_281           : integer := 281;
        s_282           : integer := 282;
        s_283           : integer := 283;
        s_284           : integer := 284;
        s_285           : integer := 285;
        s_286           : integer := 286;
        s_287           : integer := 287;
        s_288           : integer := 288;
        s_289           : integer := 289;
        s_290           : integer := 290;
        s_291           : integer := 291;
        s_292           : integer := 292;
        s_293           : integer := 293;
        s_294           : integer := 294;
        s_295           : integer := 295;
        s_296           : integer := 296;
        s_297           : integer := 297;
        s_298           : integer := 298;
        s_299           : integer := 299;
        s_300           : integer := 300;
        s_301           : integer := 301;
        s_302           : integer := 302;
        s_303           : integer := 303;
        s_304           : integer := 304;
        s_305           : integer := 305;
        s_306           : integer := 306;
        s_307           : integer := 307;
        s_308           : integer := 308;
        s_309           : integer := 309;
        s_310           : integer := 310;
        s_311           : integer := 311;
        s_312           : integer := 312;
        s_313           : integer := 313;
        s_314           : integer := 314;
        s_315           : integer := 315;
        s_316           : integer := 316;
        s_317           : integer := 317;
        s_318           : integer := 318;
        s_319           : integer := 319;
        s_320           : integer := 320;
        s_321           : integer := 321;
        s_322           : integer := 322;
        s_323           : integer := 323;
        s_324           : integer := 324;
        s_325           : integer := 325;
        s_326           : integer := 326;
        s_327           : integer := 327;
        s_328           : integer := 328;
        s_329           : integer := 329;
        s_330           : integer := 330;
        s_331           : integer := 331;
        s_332           : integer := 332;
        s_333           : integer := 333;
        s_334           : integer := 334;
        s_335           : integer := 335;
        s_336           : integer := 336;
        s_337           : integer := 337;
        s_338           : integer := 338;
        s_339           : integer := 339;
        s_340           : integer := 340;
        s_341           : integer := 341;
        s_342           : integer := 342;
        s_343           : integer := 343;
        s_344           : integer := 344;
        s_345           : integer := 345;
        s_346           : integer := 346;
        s_347           : integer := 347;
        s_348           : integer := 348;
        s_349           : integer := 349;
        s_350           : integer := 350;
        s_351           : integer := 351;
        s_352           : integer := 352;
        s_353           : integer := 353;
        s_354           : integer := 354;
        s_355           : integer := 355;
        s_356           : integer := 356;
        s_357           : integer := 357;
        s_358           : integer := 358;
        s_359           : integer := 359;
        s_360           : integer := 360;
        s_361           : integer := 361;
        s_362           : integer := 362;
        s_363           : integer := 363;
        s_364           : integer := 364;
        s_365           : integer := 365;
        s_366           : integer := 366;
        s_367           : integer := 367;
        s_368           : integer := 368;
        s_369           : integer := 369;
        s_370           : integer := 370;
        s_371           : integer := 371;
        s_372           : integer := 372;
        s_373           : integer := 373;
        s_374           : integer := 374;
        s_375           : integer := 375;
        s_376           : integer := 376;
        s_377           : integer := 377;
        s_378           : integer := 378;
        s_379           : integer := 379;
        s_380           : integer := 380;
        s_381           : integer := 381;
        s_382           : integer := 382;
        s_383           : integer := 383;
        s_384           : integer := 384;
        s_385           : integer := 385;
        s_386           : integer := 386;
        s_387           : integer := 387;
        s_388           : integer := 388;
        s_389           : integer := 389;
        s_390           : integer := 390;
        s_391           : integer := 391;
        s_392           : integer := 392;
        s_393           : integer := 393;
        s_394           : integer := 394;
        s_395           : integer := 395;
        s_396           : integer := 396;
        s_397           : integer := 397;
        s_398           : integer := 398;
        s_399           : integer := 399;
        s_400           : integer := 400;
        s_401           : integer := 401;
        s_402           : integer := 402;
        s_403           : integer := 403;
        s_404           : integer := 404;
        s_405           : integer := 405;
        s_406           : integer := 406;
        s_407           : integer := 407;
        s_408           : integer := 408;
        s_409           : integer := 409;
        s_410           : integer := 410;
        s_411           : integer := 411;
        s_412           : integer := 412;
        s_413           : integer := 413;
        s_414           : integer := 414;
        s_415           : integer := 415;
        s_416           : integer := 416;
        s_417           : integer := 417;
        s_418           : integer := 418;
        s_419           : integer := 419;
        s_420           : integer := 420;
        s_421           : integer := 421;
        s_422           : integer := 422;
        s_423           : integer := 423;
        s_424           : integer := 424;
        s_425           : integer := 425;
        s_426           : integer := 426;
        s_427           : integer := 427;
        s_428           : integer := 428;
        s_429           : integer := 429;
        s_430           : integer := 430;
        s_431           : integer := 431;
        s_432           : integer := 432;
        s_433           : integer := 433;
        s_434           : integer := 434;
        s_435           : integer := 435;
        s_436           : integer := 436;
        s_437           : integer := 437;
        s_438           : integer := 438;
        s_439           : integer := 439;
        s_440           : integer := 440;
        s_441           : integer := 441;
        s_442           : integer := 442;
        s_443           : integer := 443;
        s_444           : integer := 444;
        s_445           : integer := 445;
        s_446           : integer := 446;
        s_447           : integer := 447;
        s_448           : integer := 448;
        s_449           : integer := 449;
        s_450           : integer := 450;
        s_451           : integer := 451;
        s_452           : integer := 452;
        s_453           : integer := 453;
        s_454           : integer := 454;
        s_455           : integer := 455;
        s_456           : integer := 456;
        s_457           : integer := 457;
        s_458           : integer := 458;
        s_459           : integer := 459;
        s_460           : integer := 460;
        s_461           : integer := 461;
        s_462           : integer := 462;
        s_463           : integer := 463;
        s_464           : integer := 464;
        s_465           : integer := 465;
        s_466           : integer := 466;
        s_467           : integer := 467;
        s_468           : integer := 468;
        s_469           : integer := 469;
        s_470           : integer := 470;
        s_471           : integer := 471;
        s_472           : integer := 472;
        s_473           : integer := 473;
        s_474           : integer := 474;
        s_475           : integer := 475;
        s_476           : integer := 476;
        s_477           : integer := 477;
        s_478           : integer := 478;
        s_479           : integer := 479;
        s_480           : integer := 480;
        s_481           : integer := 481;
        s_482           : integer := 482;
        s_483           : integer := 483;
        s_484           : integer := 484;
        s_485           : integer := 485;
        s_486           : integer := 486;
        s_487           : integer := 487;
        s_488           : integer := 488;
        s_489           : integer := 489;
        s_490           : integer := 490;
        s_491           : integer := 491;
        s_492           : integer := 492;
        s_493           : integer := 493;
        s_494           : integer := 494;
        s_495           : integer := 495;
        s_496           : integer := 496;
        s_497           : integer := 497;
        s_498           : integer := 498;
        s_499           : integer := 499;
        s_500           : integer := 500;
        s_501           : integer := 501;
        s_502           : integer := 502;
        s_503           : integer := 503;
        s_504           : integer := 504;
        s_505           : integer := 505;
        s_506           : integer := 506;
        s_507           : integer := 507;
        s_508           : integer := 508;
        s_509           : integer := 509;
        s_510           : integer := 510;
        s_511           : integer := 511;
        s_512           : integer := 512;
        s_513           : integer := 513;
        s_514           : integer := 514;
        s_515           : integer := 515;
        s_516           : integer := 516;
        s_517           : integer := 517;
        s_518           : integer := 518;
        s_519           : integer := 519;
        s_520           : integer := 520;
        s_521           : integer := 521;
        s_522           : integer := 522;
        s_523           : integer := 523;
        s_524           : integer := 524;
        s_525           : integer := 525;
        s_526           : integer := 526;
        s_527           : integer := 527;
        s_528           : integer := 528;
        s_529           : integer := 529;
        s_530           : integer := 530;
        s_531           : integer := 531;
        s_532           : integer := 532;
        s_533           : integer := 533;
        s_534           : integer := 534;
        s_535           : integer := 535;
        s_536           : integer := 536;
        s_537           : integer := 537;
        s_538           : integer := 538;
        s_539           : integer := 539;
        s_540           : integer := 540;
        s_541           : integer := 541;
        s_542           : integer := 542;
        s_543           : integer := 543;
        s_544           : integer := 544;
        s_545           : integer := 545;
        s_546           : integer := 546;
        s_547           : integer := 547;
        s_548           : integer := 548;
        s_549           : integer := 549;
        s_550           : integer := 550;
        s_551           : integer := 551;
        s_552           : integer := 552;
        s_553           : integer := 553;
        s_554           : integer := 554;
        s_555           : integer := 555;
        s_556           : integer := 556;
        s_557           : integer := 557;
        s_558           : integer := 558;
        s_559           : integer := 559;
        s_560           : integer := 560;
        s_561           : integer := 561;
        s_562           : integer := 562;
        s_563           : integer := 563;
        s_564           : integer := 564;
        s_565           : integer := 565;
        s_566           : integer := 566;
        s_567           : integer := 567;
        s_568           : integer := 568;
        s_569           : integer := 569;
        s_570           : integer := 570;
        s_571           : integer := 571;
        s_572           : integer := 572;
        s_573           : integer := 573;
        s_574           : integer := 574;
        s_575           : integer := 575;
        s_576           : integer := 576;
        s_577           : integer := 577;
        s_578           : integer := 578;
        s_579           : integer := 579;
        s_580           : integer := 580;
        s_581           : integer := 581;
        s_582           : integer := 582;
        s_583           : integer := 583;
        s_584           : integer := 584;
        s_585           : integer := 585;
        s_586           : integer := 586;
        s_587           : integer := 587;
        s_588           : integer := 588;
        s_589           : integer := 589;
        s_start         : integer := 590;
        s_prefix        : integer := 591;
        s_end_error     : integer := 592;
        s_syn_error     : integer := 593
    );
    port(
        strb            : out    vl_logic;
        rw              : out    vl_logic;
        addr            : out    vl_logic_vector;
        mfc             : in     vl_logic;
        data            : inout  vl_logic_vector(7 downto 0);
        ins             : out    vl_logic_vector(2 downto 0);
        \mod\           : out    vl_logic_vector(1 downto 0);
        rm              : out    vl_logic_vector(2 downto 0);
        scale           : out    vl_logic_vector(1 downto 0);
        index_reg       : out    vl_logic_vector(2 downto 0);
        base_reg        : out    vl_logic_vector(2 downto 0);
        bits16          : out    vl_logic;
        disp            : out    vl_logic_vector;
        disp_len        : out    vl_logic_vector(2 downto 0);
        imm             : out    vl_logic_vector;
        imm_len         : out    vl_logic_vector(2 downto 0);
        bits16          : out    vl_logic;
        s               : out    vl_logic;
        w               : out    vl_logic;
        d               : out    vl_logic;
        r               : out    vl_logic;
        reg1            : out    vl_logic_vector(2 downto 0);
        reg2            : out    vl_logic_vector(2 downto 0);
        sreg2           : out    vl_logic_vector(1 downto 0);
        sreg3           : out    vl_logic_vector(2 downto 0);
        eee             : out    vl_logic_vector(2 downto 0);
        tttn            : out    vl_logic_vector(3 downto 0);
        st_i            : out    vl_logic_vector(2 downto 0);
        rdy             : out    vl_logic;
        pc_out          : out    vl_logic_vector;
        pc_in           : in     vl_logic_vector;
        reset           : in     vl_logic;
        run             : in     vl_logic;
        clk             : in     vl_logic;
        error           : out    vl_logic
    );
end idu;
